module testbench ();
   
// Declares signals for interfacing with regfile modules
    logic clock;
    logic we3;
    logic [4:0]   ra1, ra2, wa3;
    logic [31:0] rd1, rd2, wd3;
   
   integer handle3;
   integer desc3;
   logic RaR;
   
    /*logic [31:0] RefReg[31:0];
    assign RefReg[5'b00000] = 32'b00000000000000000000000000000000;
    assign RefReg[5'b00001] = 32'b00101011100101110001010010000101;
    assign RefReg[5'b00010] = 32'b00110110000111000111101001011100;
    assign RefReg[5'b00011] = 32'b10110111001010111010000011111000;
    assign RefReg[5'b00100] = 32'b11100000111111010110110001101000;
    assign RefReg[5'b00101] = 32'b01101101110001000101000010110010;
    assign RefReg[5'b00110] = 32'b00101101110011110000111110001011;
    assign RefReg[5'b00111] = 32'b11111011110101101111010001111001;
    assign RefReg[5'b01000] = 32'b11000001100011111000100001000010;
    assign RefReg[5'b01001] = 32'b01000011011010110110110011101010;
    assign RefReg[5'b01010] = 32'b00110111101000100010011011110100;
    assign RefReg[5'b01011] = 32'b01011100000111010010101111110011;
    assign RefReg[5'b01100] = 32'b00101110010100001001000011101111;
    assign RefReg[5'b01101] = 32'b01111110111001110000100000011101;
    assign RefReg[5'b01110] = 32'b11100011110010010111110010110101;
    assign RefReg[5'b01111] = 32'b11110000001110110101000101001011;
    assign RefReg[5'b10000] = 32'b00001100001111011100100100101011;
    assign RefReg[5'b10001] = 32'b00011110110100101110011110101010;
    assign RefReg[5'b10010] = 32'b01110101011010100111011010010000;
    assign RefReg[5'b10011] = 32'b10011001100110111001000110111100;
    assign RefReg[5'b10100] = 32'b11110011101011001000101000110110;
    assign RefReg[5'b10101] = 32'b10110010111011111111001001100010;
    assign RefReg[5'b10110] = 32'b10010101000010101011011110000010;
    assign RefReg[5'b10111] = 32'b00010100111000001111001000001011;
    assign RefReg[5'b11000] = 32'b01100000100101010100001101110010;
    assign RefReg[5'b11001] = 32'b01001000001100110101011011000111;
    assign RefReg[5'b11010] = 32'b00100101111110101000011110101001;
    assign RefReg[5'b11011] = 32'b00000110010110110110111011111101;
    assign RefReg[5'b11100] = 32'b10101111011100010010010110011110;
    assign RefReg[5'b11101] = 32'b11110001110110011101101000011111;
    assign RefReg[5'b11110] = 32'b10010010110011000001001111000111;
    assign RefReg[5'b11111] = 32'b10011010110010001100101000010000;

     */
   // Instantiate DUT
   regfile dut (clock,we3,ra1,ra2,wa3,wd3,rd1, rd2);

   // Setup the clock to toggle every 1 time units 
   initial 
     begin	
	clock = 1'b1;
	forever #5 clock = ~clock;
     end

   initial
     begin
	// Gives output file name
	handle3 = $fopen("rftest.out");
	// Tells when to finish simulation
	#500 $finish;		
     end

   always 
     begin
	desc3 = handle3;
	#5 $fdisplay(desc3, "%b || %b\n%b || %b\n\n", 
		   ra1, rd1, ra2, rd2);

   end   
   
   initial begin
     #0 we3 <= 1'b0; // Initialize write enable
     #0 ra1 <= 5'b0; // Initialize read addresses
     #0 ra2 <= 5'b0;
     #0 wa3 <= 5'b0; // Initialize write address
     #0 wd3 <= 420; // Initialize data to write
     
     #5 we3 <= 1'b1;
     #2 we3 <= 1'b0;
     
     #3 ra2 <= 1; // Initialize data to write
     #0 wa3 <= 1; // Initialize data to write
     #0 we3 <= 1'b1;
     #2 we3 <= 0; // Initialize data to write

/*
#5 ra1 = 5'b00000;
#0 ra2 = 5'b00000;
#0 wa3 = 5'b00000;
#0 wd3 = 32'b11111111111111111111111111111111;
#5 ra1 = 5'b00001;
#0 ra2 = 5'b00001;
#0 wa3 = 5'b00001;
#2 wd3 = 32'b00101011100101110001010010000101;
#5 ra1 = 5'b00010;
#2 ra2 = 5'b00010;
#2 wa3 = 5'b00010;
#2 wd3 = 32'b00110110000111000111101001011100;
#5 ra1 = 5'b00011;
#2 ra2 = 5'b00011;
#2 wa3 = 5'b00011;
#2 wd3 = 32'b10110111001010111010000011111000;
#5 ra1 = 5'b00100;
#2 ra2 = 5'b00100;
#2 wa3 = 5'b00100;
#2 wd3 = 32'b11100000111111010110110001101000;
#5 ra1 = 5'b00101;
#2 ra2 = 5'b00101;
#2 wa3 = 5'b00101;
#2 wd3 = 32'b01101101110001000101000010110010;
#5 ra1 = 5'b00110;
#2 ra2 = 5'b00110;
#2 wa3 = 5'b00110;
#2 wd3 = 32'b00101101110011110000111110001011;
#5 ra1 = 5'b00111;
#2 ra2 = 5'b00111;
#2 wa3 = 5'b00111;
#2 wd3 = 32'b11111011110101101111010001111001;
#5 ra1 = 5'b01000;
#2 ra2 = 5'b01000;
#2 wa3 = 5'b01000;
#2 wd3 = 32'b11000001100011111000100001000010;
#5 ra1 = 5'b01001;
#2 ra2 = 5'b01001;
#2 wa3 = 5'b01001;
#2 wd3 = 32'b01000011011010110110110011101010;
#5 ra1 = 5'b01010;
#2 ra2 = 5'b01010;
#2 wa3 = 5'b01010;
#2 wd3 = 32'b00110111101000100010011011110100;
#5 ra1 = 5'b01011;
#2 ra2 = 5'b01011;
#2 wa3 = 5'b01011;
#2 wd3 = 32'b01011100000111010010101111110011;
#5 ra1 = 5'b01100;
#2 ra2 = 5'b01100;
#2 wa3 = 5'b01100;
#2 wd3 = 32'b00101110010100001001000011101111;
#5 ra1 = 5'b01101;
#2 ra2 = 5'b01101;
#2 wa3 = 5'b01101;
#2 wd3 = 32'b01111110111001110000100000011101;
#5 ra1 = 5'b01110;
#2 ra2 = 5'b01110;
#2 wa3 = 5'b01110;
#2 wd3 = 32'b11100011110010010111110010110101;
#5 ra1 = 5'b01111;
#2 ra2 = 5'b01111;
#2 wa3 = 5'b01111;
#2 wd3 = 32'b11110000001110110101000101001011;
#5 ra1 = 5'b10000;
#2 ra2 = 5'b10000;
#2 wa3 = 5'b10000;
#2 wd3 = 32'b00001100001111011100100100101011;
#5 ra1 = 5'b10001;
#2 ra2 = 5'b10001;
#2 wa3 = 5'b10001;
#2 wd3 = 32'b00011110110100101110011110101010;
#5 ra1 = 5'b10010;
#2 ra2 = 5'b10010;
#2 wa3 = 5'b10010;
#2 wd3 = 32'b01110101011010100111011010010000;
#5 ra1 = 5'b10011;
#2 ra2 = 5'b10011;
#2 wa3 = 5'b10011;
#2 wd3 = 32'b10011001100110111001000110111100;
#5 ra1 = 5'b10100;
#2 ra2 = 5'b10100;
#2 wa3 = 5'b10100;
#2 wd3 = 32'b11110011101011001000101000110110;
#5 ra1 = 5'b10101;
#2 ra2 = 5'b10101;
#2 wa3 = 5'b10101;
#2 wd3 = 32'b10110010111011111111001001100010;
#5 ra1 = 5'b10110;
#2 ra2 = 5'b10110;
#2 wa3 = 5'b10110;
#2 wd3 = 32'b10010101000010101011011110000010;
#5 ra1 = 5'b10111;
#2 ra2 = 5'b10111;
#2 wa3 = 5'b10111;
#2 wd3 = 32'b00010100111000001111001000001011;
#5 ra1 = 5'b11000;
#2 ra2 = 5'b11000;
#2 wa3 = 5'b11000;
#2 wd3 = 32'b01100000100101010100001101110010;
#5 ra1 = 5'b11001;
#2 ra2 = 5'b11001;
#2 wa3 = 5'b11001;
#2 wd3 = 32'b01001000001100110101011011000111;
#5 ra1 = 5'b11010;
#2 ra2 = 5'b11010;
#2 wa3 = 5'b11010;
#2 wd3 = 32'b00100101111110101000011110101001;
#5 ra1 = 5'b11011;
#2 ra2 = 5'b11011;
#2 wa3 = 5'b11011;
#2 wd3 = 32'b00000110010110110110111011111101;
#5 ra1 = 5'b11100;
#2 ra2 = 5'b11100;
#2 wa3 = 5'b11100;
#2 wd3 = 32'b10101111011100010010010110011110;
#5 ra1 = 5'b11101;
#2 ra2 = 5'b11101;
#2 wa3 = 5'b11101;
#2 wd3 = 32'b11110001110110011101101000011111;
#5 ra1 = 5'b11110;
#2 ra2 = 5'b11110;
#2 wa3 = 5'b11110;
#2 wd3 = 32'b10010010110011000001001111000111;
#5 ra1 = 5'b11111;
#2 ra2 = 5'b11111;
#2 wa3 = 5'b11111;
#2 wd3 = 32'b10011010110010001100101000010000;


/*
     #5 ra1, ra2, wa3 = 5'b00001;
     #5 wd3 = 32'b00101011100101110001010010000101;
     #5 ra1, ra2, wa3 = 5'b00010;
     #5 wd3 = 32'b00110110000111000111101001011100;
     #5 ra1, ra2, wa3 = 5'b00011;
     #5 wd3 = 32'b10110111001010111010000011111000;
     #5 ra1, ra2, wa3 = 5'b00100;
     #5 wd3 = 32'b11100000111111010110110001101000;
     #5 ra1, ra2, wa3 = 5'b00101;
     #5 wd3 = 32'b01101101110001000101000010110010;
     #5 ra1, ra2, wa3 = 5'b00110;
     #5 wd3 = 32'b00101101110011110000111110001011;
     #5 ra1, ra2, wa3 = 5'b00111;
     #5 wd3 = 32'b11111011110101101111010001111001;
     #5 ra1, ra2, wa3 = 5'b01000;
     #5 wd3 = 32'b11000001100011111000100001000010;
     #5 ra1, ra2, wa3 = 5'b01001;
     #5 wd3 = 32'b01000011011010110110110011101010;
     #5 ra1, ra2, wa3 = 5'b01010;
     #5 wd3 = 32'b00110111101000100010011011110100;
     #5 ra1, ra2, wa3 = 5'b01011;
     #5 wd3 = 32'b01011100000111010010101111110011;
     #5 ra1, ra2, wa3 = 5'b01100;
     #5 wd3 = 32'b00101110010100001001000011101111;
     #5 ra1, ra2, wa3 = 5'b01101;
     #5 wd3 = 32'b01111110111001110000100000011101;
     #5 ra1, ra2, wa3 = 5'b01110;
     #5 wd3 = 32'b11100011110010010111110010110101;
     #5 ra1, ra2, wa3 = 5'b01111;
     #5 wd3 = 32'b11110000001110110101000101001011;
     #5 ra1, ra2, wa3 = 5'b10000;
     #5 wd3 = 32'b00001100001111011100100100101011;
     #5 ra1, ra2, wa3 = 5'b10001;
     #5 wd3 = 32'b00011110110100101110011110101010;
     #5 ra1, ra2, wa3 = 5'b10010;
     #5 wd3 = 32'b01110101011010100111011010010000;
     #5 ra1, ra2, wa3 = 5'b10011;
     #5 wd3 = 32'b10011001100110111001000110111100;
     #5 ra1, ra2, wa3 = 5'b10100;
     #5 wd3 = 32'b11110011101011001000101000110110;
     #5 ra1, ra2, wa3 = 5'b10101;
     #5 wd3 = 32'b10110010111011111111001001100010;
     #5 ra1, ra2, wa3 = 5'b10110;
     #5 wd3 = 32'b10010101000010101011011110000010;
     #5 ra1, ra2, wa3 = 5'b10111;
     #5 wd3 = 32'b00010100111000001111001000001011;
     #5 ra1, ra2, wa3 = 5'b11000;
     #5 wd3 = 32'b01100000100101010100001101110010;
     #5 ra1, ra2, wa3 = 5'b11001;
     #5 wd3 = 32'b01001000001100110101011011000111;
     #5 ra1, ra2, wa3 = 5'b11010;
     #5 wd3 = 32'b00100101111110101000011110101001;
     #5 ra1, ra2, wa3 = 5'b11011;
     #5 wd3 = 32'b00000110010110110110111011111101;
     #5 ra1, ra2, wa3 = 5'b11100;
     #5 wd3 = 32'b10101111011100010010010110011110;
     #5 ra1, ra2, wa3 = 5'b11101;
     #5 wd3 = 32'b11110001110110011101101000011111;
     #5 ra1, ra2, wa3 = 5'b11110;
     #5 wd3 = 32'b10010010110011000001001111000111;
     #5 ra1, ra2, wa3 = 5'b11111;
     #5 wd3 = 32'b10011010110010001100101000010000;
     /*#5 ra1 = 5'b00000;
     #5 ra1 = 5'b00001;
     #5 ra1 = 5'b00010;
     #5 ra1 = 5'b00011;
     #5 ra1 = 5'b00100;
     #5 ra1 = 5'b00101;
     #5 ra1 = 5'b00110;
     #5 ra1 = 5'b00111;
     #5 ra1 = 5'b01000;
     #5 ra1 = 5'b01001;
     #5 ra1 = 5'b01010;
     #5 ra1 = 5'b01011;
     #5 ra1 = 5'b01100;
     #5 ra1 = 5'b01101;
     #5 ra1 = 5'b01110;
     #5 ra1 = 5'b01111;
     #5 ra1 = 5'b10000;
     #5 ra1 = 5'b10001;
     #5 ra1 = 5'b10010;
     #5 ra1 = 5'b10011;
     #5 ra1 = 5'b10100;
     #5 ra1 = 5'b10101;
     #5 ra1 = 5'b10110;
     #5 ra1 = 5'b10111;
     #5 ra1 = 5'b11000;
     #5 ra1 = 5'b11001;
     #5 ra1 = 5'b11010;
     #5 ra1 = 5'b11011;
     #5 ra1 = 5'b11100;
     #5 ra1 = 5'b11101;
     #5 ra1 = 5'b11110;

     #5 ra1 = 5'b11111;  
     #5 ra2 = 5'b00000;
     #5 ra2 = 5'b00001;
     #5 ra2 = 5'b00010;
     #5 ra2 = 5'b00011;
     #5 ra2 = 5'b00100;
     #5 ra2 = 5'b00101;
     #5 ra2 = 5'b00110;
     #5 ra2 = 5'b00111;
     #5 ra2 = 5'b01000;
     #5 ra2 = 5'b01001;
     #5 ra2 = 5'b01010;
     #5 ra2 = 5'b01011;
     #5 ra2 = 5'b01100;
     #5 ra2 = 5'b01101;
     #5 ra2 = 5'b01110;
     #5 ra2 = 5'b01111;
     #5 ra2 = 5'b10000;
     #5 ra2 = 5'b10001;
     #5 ra2 = 5'b10010;
     #5 ra2 = 5'b10011;
     #5 ra2 = 5'b10100;
     #5 ra2 = 5'b10101;
     #5 ra2 = 5'b10110;
     #5 ra2 = 5'b10111;
     #5 ra2 = 5'b11000;
     #5 ra2 = 5'b11001;
     #5 ra2 = 5'b11010;
     #5 ra2 = 5'b11011;
     #5 ra2 = 5'b11100;
     #5 ra2 = 5'b11101;
     #5 ra2 = 5'b11110;
     #5 ra2 = 5'b11111;
     */
     #3 we3 = 1'b0; // Set write enable low
     
      // Write data to register file
     //for (i = 0; i < 32; i = i+) begin
     //    #2 wa3 = i;
     //    #2 wd3 = 69;
     //    #2;
     // end


      // Read data from register file
     //for (i = 0; i < 32; i++) begin
     //    #1 ra1 = i;
     //    #1; // You may need a delay here to observe the output
     //end
     




   end

endmodule // regfile

